module comparator(a1,a2,b1,b2,y1,y2);//???? ??

input[2:0] a1,a2,b1,b2;//3bit input a1,a2,b1,b2
output y1,y2;//output y1,y2
reg y1,y2;//register value y1,y2

always@(a1 or a2 or b1 or b2)//a1,a2,b1,b2 ? ?? ??? ?? ??? ?? ??

begin

if(a1[0]==a2[0])//0? ?? ??, ?? ?? else ? ?? y1=0(L17)
	if(a1[1]==a2[1])//1? ?? ??, ?? ?? else ? ?? y1=0(L16)
		if(a1[2]==a2[2])//2? ?? ??, ?? ?? y1=1 ?? ?? else ? ?? y1=0(L15)
			y1=1;
else y1=0;

if(b1==b2)//b1,b2? ??
	y2=1;
else
	y2=0;//??? y2=1, ??? y2=0
end 
endmodule