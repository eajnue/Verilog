module evenparity(a,z);//????
 
input[7:0] a;//8bit intput a
output[8:0] z;//9bit output z
reg[8:0] z;//9bit reg vaue z

always@(a)//a? ?? ??? ??
begin

z[8:1]<=a[7:0];//z? 1?~8? ??? a? 0?~7? ??? ? ??

if(^a[7:0]) z[0]<=1;//a?? 1? ??? ???? z? 0? ?? 1
else z[0]<=0;//a?? 1? ??? ???? z? 0? ?? 0 

end

endmodule




















































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































