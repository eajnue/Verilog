module and_module(a,b,z);

input a,b;
output z;

wire z;

and a1(z,a,b);

endmodule

